`include "uart_trx.v"

//----------------------------------------------------------------------------
//                                                                          --
//                         Module Declaration                               --
//                                                                          --
//----------------------------------------------------------------------------
module top (
  // outputs
  //output wire led_red  , 
  // Red
  //output wire led_blue , 
  // Blue
  //output wire led_green , 
  // Green
  output wire uarttx , 
  // UART Transmission pin
  //input wire uartrx , 
  // UART Transmission pin
  input wire  hw_clk,
  input  wire sensor_in
);

  //wire        int_osc            ;
  //reg  [27:0] frequency_counter_i;
  
/* 9600 Hz clock generation (from 12 MHz) */
    reg clk_9600 = 0;
    reg [31:0] divcnt = 0;
    //reg [31:0] cntr_9600 = 32'b0;
    localparam DIV = 625;
    //parameter period_9600 = 625;
    
//uart_tx_8n1 DanUART (.clk (clk_9600), .txbyte("D"), .senddata(frequency_counter_i[24]), .tx(uarttx));
//----------------------------------------------------------------------------
//                                                                          --
//                       Internal Oscillator                                --
//                                                                          --
//----------------------------------------------------------------------------
  //SB_HFOSC #(.CLKHF_DIV ("0b10")) u_SB_HFOSC ( .CLKHFPU(1'b1), .CLKHFEN(1'b1), .CLKHF(int_osc));


//----------------------------------------------------------------------------
//                                                                          --
//                       Counter                                            --
//                                                                          --
//----------------------------------------------------------------------------

always @(posedge hw_clk) begin
    if (divcnt == DIV) begin
      clk_9600 <= ~clk_9600;
      divcnt    <= 0;
    end else
      divcnt <= divcnt + 1;
  end

  //always @(posedge int_osc) begin
    //frequency_counter_i <= frequency_counter_i + 1'b1;
        /* generate 9600 Hz clock */
        //cntr_9600 <= cntr_9600 + 1;
        //if (cntr_9600 == period_9600) begin
            //clk_9600 <= ~clk_9600;
            //cntr_9600 <= 32'b0;
        //end
  //end

reg prev_sample = 1;
  reg send_pulse  = 0;
  always @(posedge clk_9600) begin
    if (sensor_in != prev_sample) begin
      send_pulse  <= 1;
      prev_sample <= sensor_in;
    end else
      send_pulse <= 0;
  end

wire [7:0] txbyte = (prev_sample) ? "1" : "0";

//----------------------------------------------------------------------------
//                                                                          --
//                       Instantiate RGB primitive                          --
//                                                                          --
//----------------------------------------------------------------------------
  //SB_RGBA_DRV RGB_DRIVER (
    //.RGBLEDEN(1'b1                                            ),
    //.RGB0PWM (uartrx),
    //.RGB1PWM (uartrx),
    //.RGB2PWM (uartrx),
    //.CURREN  (1'b1                                            ),
    //.RGB0    (led_green                                       ), 
//Actual Hardware connection
    //.RGB1    (led_blue                                        ),
    //.RGB2    (led_red                                         )
  //);
  //defparam RGB_DRIVER.RGB0_CURRENT = "0b000001";
  //defparam RGB_DRIVER.RGB1_CURRENT = "0b000001";
  //defparam RGB_DRIVER.RGB2_CURRENT = "0b000001";

 uart_tx_8n1 U1 (
    .clk      (clk_9600),
    .txbyte   (txbyte),
    .senddata (send_pulse),
    .tx       (uarttx)
  );

endmodule
