//`include "uart_trx.v"

//----------------------------------------------------------------------------
//                                                                          --
//                         Module Declaration                               --
//                                                                          --
//----------------------------------------------------------------------------
module top (
  // outputs
  output wire led_red  , // Red
  output wire led_blue , // Blue
  output wire led_green , // Green
  output wire uarttx , // UART Transmission pin
  input wire  hw_clk
);

  //wire        int_osc            ;
  wire clk_main = hw_clk;
  reg  [27:0] frequency_counter_i;
  
/* 9600 Hz clock generation (from 12 MHz) */
    reg clk_9600 = 0;
    reg [31:0] cntr_9600 = 32'b0;
    parameter period_9600 = 625;
    
uart_tx_8n1 DanUART (.clk (clk_9600), .txbyte("D"), .senddata(frequency_counter_i[24]), .tx(uarttx));
//----------------------------------------------------------------------------
//                                                                          --
//                       Internal Oscillator                                --
//                                                                          --
//----------------------------------------------------------------------------
  //SB_HFOSC #(.CLKHF_DIV ("0b10")) u_SB_HFOSC //( .CLKHFPU(1'b1), .CLKHFEN(1'b1), .CLKHF(int_osc));


//----------------------------------------------------------------------------
//                                                                          --
//                       Counter                                            --
//                                                                          --
//----------------------------------------------------------------------------
  //always @(posedge int_osc) begin
  always @(posedge clk_main) begin
    frequency_counter_i <= frequency_counter_i + 1'b1;
        /* generate 9600 Hz clock */
        cntr_9600 <= cntr_9600 + 1;
        if (cntr_9600 == period_9600) begin
            clk_9600 <= ~clk_9600;
            cntr_9600 <= 32'b0;
        end
  end

//----------------------------------------------------------------------------
//                                                                          --
//                       Instantiate RGB primitive                          --
//                                                                          --
//----------------------------------------------------------------------------
  //SB_RGBA_DRV RGB_DRIVER (
  //  .RGBLEDEN(1'b1                                            ),
  //  .RGB0PWM (frequency_counter_i[24]&frequency_counter_i[23] ),
  //  .RGB1PWM (frequency_counter_i[24]&~frequency_counter_i[23]),
  //  .RGB2PWM (~frequency_counter_i[24]&frequency_counter_i[23]),
  //  .CURREN  (1'b1                                            ),
  //  .RGB0    (led_green                                       ), 
  //Actual Hardware connection
  //  .RGB1    (led_blue                                        ),
  //  .RGB2    (led_red                                         )
  //);
  //defparam RGB_DRIVER.RGB0_CURRENT = "0b000001";
  //defparam RGB_DRIVER.RGB1_CURRENT = "0b000001";
  //defparam RGB_DRIVER.RGB2_CURRENT = "0b000001";

  assign led_green = frequency_counter_i[24] & frequency_counter_i[23];
  assign led_blue  = frequency_counter_i[24] & ~frequency_counter_i[23];
  assign led_red   = ~frequency_counter_i[24] & frequency_counter_i[23];

endmodule
